* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colend.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colend BL1 VPWR VGND BL0
X0 BL0 a_0_24# BL0 VGND sky130_fd_pr__special_nfet_pass w=0.07u l=0.21u
.ends
