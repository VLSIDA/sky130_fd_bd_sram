* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colenda.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colenda bl vdd gnd br gate vpb vnb
X0 br gate br vnb sky130_fd_pr__special_nfet_pass w=0.065u l=0.17u
.ends

