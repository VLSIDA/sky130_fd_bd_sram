* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colend.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_colend_replica bl br vdd gnd vpb vnb gate
X0 br gate br vnb sky130_fd_pr__special_nfet_pass w=0.14u l=0.14u
.ends
