* NGSPICE file created from sky130_fd_bd_sram__openram_sp_cell_opt1_dummy.ext - technology: sky130A
.subckt sky130_fd_bd_sram__openram_sp_cell_opt1_dummy BL BR VGND VPWR VPB VNB WL

*inverter 1
X6 Q Q_bar VPWR VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X1 Q Q_bar VGND VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15

*inverter 2
X5 VPWR Q Q_bar VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X7 VGND Q Q_bar VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15

*access tx
X2 Q wl bl_noconn VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
X0 Q_bar wl br_noconn VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15

X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass w=0.14 l=25n
X4 Q_bar WL Q_bar VPB sky130_fd_pr__special_pfet_pass w=0.14 l=25n
.ends
