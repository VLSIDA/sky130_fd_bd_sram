* NGSPICE file created from sky130_fd_bd_sram__openram_sp_cell_opt1_dummy.ext - technology: sky130A
.subckt sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy BL BR VGND VPWR VPB VNB WL

*inverter 1
X6 VPWR VGND lr_parasitic_float VPB sky130_fd_pr__special_pfet_pass w=0.14u l=0.15u
X1 VGND VGND ll_access_float VNB sky130_fd_pr__special_nfet_latch w=0.21u l=0.15u

*inverter 2
X5 VPWR VGND ur_parasitic_float VPB sky130_fd_pr__special_pfet_pass w=0.14u l=0.15u
X7 VGND VGND ul_access_float VNB sky130_fd_pr__special_nfet_latch w=0.21u l=0.15u

*access tx
X2 ul_access_float WL BL VNB sky130_fd_pr__special_nfet_pass w=0.14u l=0.15u
X0 ll_access_float WL BR VNB sky130_fd_pr__special_nfet_pass w=0.14u l=0.15u

X3 ur_parasitic_float WL ur_parasitic_float VPB sky130_fd_pr__special_pfet_pass w=0.14u l=25n
X4 lr_parasitic_float WL lr_parasitic_float VPB sky130_fd_pr__special_pfet_pass w=0.14u l=25n
.ends
