* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* NGSPICE file created from sky130_fd_bd_sram__openram_sp_nand4_dec.ext - technology: EFS8A

.subckt sky130_fd_bd_sram__openram_sp_nand4_dec A B C D Z VDD GND
M1000 Z A a_406_334# GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15 m=1 mult=1
M1004 a_406_190# D GND GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15 m=1 mult=1
M1005 a_406_262# C a_406_190# GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15 m=1 mult=1
M1007 a_406_334# B a_406_262# GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15 m=1 mult=1
M1001 Z A VDD VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15 m=1 mult=1
M1002 VDD C Z VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15 m=1 mult=1
M1003 VDD D Z VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15 m=1 mult=1
M1006 Z B VDD VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15 m=1 mult=1
.ends

