* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Ingore first line
.SUBCKT sky130_fd_bd_sram__openram_dp_cell_replica BL0 BR0 BL1 BR1 WL0 WL1 VDD GND
** N=9 EP=8 IP=0 FDC=16
*.SEEDPROM

* Bitcell Core
M0 Q WL1 BL1 GND sky130_fd_pr__nfet_01v8 W=0.21u L=0.15u m=1 mult=1
M1 GND VDD Q GND sky130_fd_pr__nfet_01v8 W=0.21u L=0.15u m=1 mult=1
M2 GND VDD Q GND sky130_fd_pr__nfet_01v8 W=0.21u L=0.15u m=1 mult=1
M3 BL0 WL0 Q GND sky130_fd_pr__nfet_01v8 W=0.21u L=0.15u m=1 mult=1
M4 VDD WL1 BR1 GND sky130_fd_pr__nfet_01v8 W=0.21u L=0.15u m=1 mult=1
M5 GND Q VDD GND sky130_fd_pr__nfet_01v8 W=0.21u L=0.15u m=1 mult=1
M6 GND Q VDD GND sky130_fd_pr__nfet_01v8 W=0.21u L=0.15u m=1 mult=1
M7 BR0 WL0 VDD GND sky130_fd_pr__nfet_01v8 W=0.21u L=0.15u m=1 mult=1
M8 VDD Q VDD VDD sky130_fd_pr__pfet_01v8_hvt W=0.14u L=0.15u m=1 mult=1
M9 Q VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt W=0.14u L=0.15u m=1 mult=1

* drainOnly PMOS
*M10 VDD WL1 VDD VDD sky130_fd_pr__pfet_01v8_hvtu L=0.08 W=0.14u m=1 mult=1
*M11 Q WL0 Q VDD sky130_fd_pr__pfet_01v8_hvtu L=0.08 W=0.14u m=1 mult=1

* drainOnly NMOS
*M12 BL1 GND BL1 GND sky130_fd_pr__nfet_01v8 W=0.21u L=0.08u m=1 mult=1
*M14 BR1 GND BR1 GND sky130_fd_pr__nfet_01v8 W=0.21u L=0.08u m=1 mult=1

.ENDS
